magic
tech sky130A
magscale 1 2
timestamp 1716975249
<< obsli1 >>
rect 1104 2159 438840 437393
<< obsm1 >>
rect 934 1368 438840 437424
<< metal2 >>
rect 16210 0 16266 800
rect 17038 0 17094 800
rect 17866 0 17922 800
rect 18694 0 18750 800
rect 19522 0 19578 800
rect 20350 0 20406 800
rect 21178 0 21234 800
rect 22006 0 22062 800
rect 22834 0 22890 800
rect 23662 0 23718 800
rect 24490 0 24546 800
rect 25318 0 25374 800
rect 26146 0 26202 800
rect 26974 0 27030 800
rect 27802 0 27858 800
rect 28630 0 28686 800
rect 29458 0 29514 800
rect 30286 0 30342 800
rect 31114 0 31170 800
rect 31942 0 31998 800
rect 32770 0 32826 800
rect 33598 0 33654 800
rect 34426 0 34482 800
rect 35254 0 35310 800
rect 36082 0 36138 800
rect 36910 0 36966 800
rect 37738 0 37794 800
rect 38566 0 38622 800
rect 39394 0 39450 800
rect 40222 0 40278 800
rect 41050 0 41106 800
rect 41878 0 41934 800
rect 42706 0 42762 800
rect 43534 0 43590 800
rect 44362 0 44418 800
rect 45190 0 45246 800
rect 46018 0 46074 800
rect 46846 0 46902 800
rect 47674 0 47730 800
rect 48502 0 48558 800
rect 49330 0 49386 800
rect 50158 0 50214 800
rect 50986 0 51042 800
rect 51814 0 51870 800
rect 52642 0 52698 800
rect 53470 0 53526 800
rect 54298 0 54354 800
rect 55126 0 55182 800
rect 55954 0 56010 800
rect 56782 0 56838 800
rect 57610 0 57666 800
rect 58438 0 58494 800
rect 59266 0 59322 800
rect 60094 0 60150 800
rect 60922 0 60978 800
rect 61750 0 61806 800
rect 62578 0 62634 800
rect 63406 0 63462 800
rect 64234 0 64290 800
rect 65062 0 65118 800
rect 65890 0 65946 800
rect 66718 0 66774 800
rect 67546 0 67602 800
rect 68374 0 68430 800
rect 69202 0 69258 800
rect 70030 0 70086 800
rect 70858 0 70914 800
rect 71686 0 71742 800
rect 72514 0 72570 800
rect 73342 0 73398 800
rect 74170 0 74226 800
rect 74998 0 75054 800
rect 75826 0 75882 800
rect 76654 0 76710 800
rect 77482 0 77538 800
rect 78310 0 78366 800
rect 79138 0 79194 800
rect 79966 0 80022 800
rect 80794 0 80850 800
rect 81622 0 81678 800
rect 82450 0 82506 800
rect 83278 0 83334 800
rect 84106 0 84162 800
rect 84934 0 84990 800
rect 85762 0 85818 800
rect 86590 0 86646 800
rect 87418 0 87474 800
rect 88246 0 88302 800
rect 89074 0 89130 800
rect 89902 0 89958 800
rect 90730 0 90786 800
rect 91558 0 91614 800
rect 92386 0 92442 800
rect 93214 0 93270 800
rect 94042 0 94098 800
rect 94870 0 94926 800
rect 95698 0 95754 800
rect 96526 0 96582 800
rect 97354 0 97410 800
rect 98182 0 98238 800
rect 99010 0 99066 800
rect 99838 0 99894 800
rect 100666 0 100722 800
rect 101494 0 101550 800
rect 102322 0 102378 800
rect 103150 0 103206 800
rect 103978 0 104034 800
rect 104806 0 104862 800
rect 105634 0 105690 800
rect 106462 0 106518 800
rect 107290 0 107346 800
rect 108118 0 108174 800
rect 108946 0 109002 800
rect 109774 0 109830 800
rect 110602 0 110658 800
rect 111430 0 111486 800
rect 112258 0 112314 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115570 0 115626 800
rect 116398 0 116454 800
rect 117226 0 117282 800
rect 118054 0 118110 800
rect 118882 0 118938 800
rect 119710 0 119766 800
rect 120538 0 120594 800
rect 121366 0 121422 800
rect 122194 0 122250 800
rect 123022 0 123078 800
rect 123850 0 123906 800
rect 124678 0 124734 800
rect 125506 0 125562 800
rect 126334 0 126390 800
rect 127162 0 127218 800
rect 127990 0 128046 800
rect 128818 0 128874 800
rect 129646 0 129702 800
rect 130474 0 130530 800
rect 131302 0 131358 800
rect 132130 0 132186 800
rect 132958 0 133014 800
rect 133786 0 133842 800
rect 134614 0 134670 800
rect 135442 0 135498 800
rect 136270 0 136326 800
rect 137098 0 137154 800
rect 137926 0 137982 800
rect 138754 0 138810 800
rect 139582 0 139638 800
rect 140410 0 140466 800
rect 141238 0 141294 800
rect 142066 0 142122 800
rect 142894 0 142950 800
rect 143722 0 143778 800
rect 144550 0 144606 800
rect 145378 0 145434 800
rect 146206 0 146262 800
rect 147034 0 147090 800
rect 147862 0 147918 800
rect 148690 0 148746 800
rect 149518 0 149574 800
rect 150346 0 150402 800
rect 151174 0 151230 800
rect 152002 0 152058 800
rect 152830 0 152886 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155314 0 155370 800
rect 156142 0 156198 800
rect 156970 0 157026 800
rect 157798 0 157854 800
rect 158626 0 158682 800
rect 159454 0 159510 800
rect 160282 0 160338 800
rect 161110 0 161166 800
rect 161938 0 161994 800
rect 162766 0 162822 800
rect 163594 0 163650 800
rect 164422 0 164478 800
rect 165250 0 165306 800
rect 166078 0 166134 800
rect 166906 0 166962 800
rect 167734 0 167790 800
rect 168562 0 168618 800
rect 169390 0 169446 800
rect 170218 0 170274 800
rect 171046 0 171102 800
rect 171874 0 171930 800
rect 172702 0 172758 800
rect 173530 0 173586 800
rect 174358 0 174414 800
rect 175186 0 175242 800
rect 176014 0 176070 800
rect 176842 0 176898 800
rect 177670 0 177726 800
rect 178498 0 178554 800
rect 179326 0 179382 800
rect 180154 0 180210 800
rect 180982 0 181038 800
rect 181810 0 181866 800
rect 182638 0 182694 800
rect 183466 0 183522 800
rect 184294 0 184350 800
rect 185122 0 185178 800
rect 185950 0 186006 800
rect 186778 0 186834 800
rect 187606 0 187662 800
rect 188434 0 188490 800
rect 189262 0 189318 800
rect 190090 0 190146 800
rect 190918 0 190974 800
rect 191746 0 191802 800
rect 192574 0 192630 800
rect 193402 0 193458 800
rect 194230 0 194286 800
rect 195058 0 195114 800
rect 195886 0 195942 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198370 0 198426 800
rect 199198 0 199254 800
rect 200026 0 200082 800
rect 200854 0 200910 800
rect 201682 0 201738 800
rect 202510 0 202566 800
rect 203338 0 203394 800
rect 204166 0 204222 800
rect 204994 0 205050 800
rect 205822 0 205878 800
rect 206650 0 206706 800
rect 207478 0 207534 800
rect 208306 0 208362 800
rect 209134 0 209190 800
rect 209962 0 210018 800
rect 210790 0 210846 800
rect 211618 0 211674 800
rect 212446 0 212502 800
rect 213274 0 213330 800
rect 214102 0 214158 800
rect 214930 0 214986 800
rect 215758 0 215814 800
rect 216586 0 216642 800
rect 217414 0 217470 800
rect 218242 0 218298 800
rect 219070 0 219126 800
rect 219898 0 219954 800
rect 220726 0 220782 800
rect 221554 0 221610 800
rect 222382 0 222438 800
rect 223210 0 223266 800
rect 224038 0 224094 800
rect 224866 0 224922 800
rect 225694 0 225750 800
rect 226522 0 226578 800
rect 227350 0 227406 800
rect 228178 0 228234 800
rect 229006 0 229062 800
rect 229834 0 229890 800
rect 230662 0 230718 800
rect 231490 0 231546 800
rect 232318 0 232374 800
rect 233146 0 233202 800
rect 233974 0 234030 800
rect 234802 0 234858 800
rect 235630 0 235686 800
rect 236458 0 236514 800
rect 237286 0 237342 800
rect 238114 0 238170 800
rect 238942 0 238998 800
rect 239770 0 239826 800
rect 240598 0 240654 800
rect 241426 0 241482 800
rect 242254 0 242310 800
rect 243082 0 243138 800
rect 243910 0 243966 800
rect 244738 0 244794 800
rect 245566 0 245622 800
rect 246394 0 246450 800
rect 247222 0 247278 800
rect 248050 0 248106 800
rect 248878 0 248934 800
rect 249706 0 249762 800
rect 250534 0 250590 800
rect 251362 0 251418 800
rect 252190 0 252246 800
rect 253018 0 253074 800
rect 253846 0 253902 800
rect 254674 0 254730 800
rect 255502 0 255558 800
rect 256330 0 256386 800
rect 257158 0 257214 800
rect 257986 0 258042 800
rect 258814 0 258870 800
rect 259642 0 259698 800
rect 260470 0 260526 800
rect 261298 0 261354 800
rect 262126 0 262182 800
rect 262954 0 263010 800
rect 263782 0 263838 800
rect 264610 0 264666 800
rect 265438 0 265494 800
rect 266266 0 266322 800
rect 267094 0 267150 800
rect 267922 0 267978 800
rect 268750 0 268806 800
rect 269578 0 269634 800
rect 270406 0 270462 800
rect 271234 0 271290 800
rect 272062 0 272118 800
rect 272890 0 272946 800
rect 273718 0 273774 800
rect 274546 0 274602 800
rect 275374 0 275430 800
rect 276202 0 276258 800
rect 277030 0 277086 800
rect 277858 0 277914 800
rect 278686 0 278742 800
rect 279514 0 279570 800
rect 280342 0 280398 800
rect 281170 0 281226 800
rect 281998 0 282054 800
rect 282826 0 282882 800
rect 283654 0 283710 800
rect 284482 0 284538 800
rect 285310 0 285366 800
rect 286138 0 286194 800
rect 286966 0 287022 800
rect 287794 0 287850 800
rect 288622 0 288678 800
rect 289450 0 289506 800
rect 290278 0 290334 800
rect 291106 0 291162 800
rect 291934 0 291990 800
rect 292762 0 292818 800
rect 293590 0 293646 800
rect 294418 0 294474 800
rect 295246 0 295302 800
rect 296074 0 296130 800
rect 296902 0 296958 800
rect 297730 0 297786 800
rect 298558 0 298614 800
rect 299386 0 299442 800
rect 300214 0 300270 800
rect 301042 0 301098 800
rect 301870 0 301926 800
rect 302698 0 302754 800
rect 303526 0 303582 800
rect 304354 0 304410 800
rect 305182 0 305238 800
rect 306010 0 306066 800
rect 306838 0 306894 800
rect 307666 0 307722 800
rect 308494 0 308550 800
rect 309322 0 309378 800
rect 310150 0 310206 800
rect 310978 0 311034 800
rect 311806 0 311862 800
rect 312634 0 312690 800
rect 313462 0 313518 800
rect 314290 0 314346 800
rect 315118 0 315174 800
rect 315946 0 316002 800
rect 316774 0 316830 800
rect 317602 0 317658 800
rect 318430 0 318486 800
rect 319258 0 319314 800
rect 320086 0 320142 800
rect 320914 0 320970 800
rect 321742 0 321798 800
rect 322570 0 322626 800
rect 323398 0 323454 800
rect 324226 0 324282 800
rect 325054 0 325110 800
rect 325882 0 325938 800
rect 326710 0 326766 800
rect 327538 0 327594 800
rect 328366 0 328422 800
rect 329194 0 329250 800
rect 330022 0 330078 800
rect 330850 0 330906 800
rect 331678 0 331734 800
rect 332506 0 332562 800
rect 333334 0 333390 800
rect 334162 0 334218 800
rect 334990 0 335046 800
rect 335818 0 335874 800
rect 336646 0 336702 800
rect 337474 0 337530 800
rect 338302 0 338358 800
rect 339130 0 339186 800
rect 339958 0 340014 800
rect 340786 0 340842 800
rect 341614 0 341670 800
rect 342442 0 342498 800
rect 343270 0 343326 800
rect 344098 0 344154 800
rect 344926 0 344982 800
rect 345754 0 345810 800
rect 346582 0 346638 800
rect 347410 0 347466 800
rect 348238 0 348294 800
rect 349066 0 349122 800
rect 349894 0 349950 800
rect 350722 0 350778 800
rect 351550 0 351606 800
rect 352378 0 352434 800
rect 353206 0 353262 800
rect 354034 0 354090 800
rect 354862 0 354918 800
rect 355690 0 355746 800
rect 356518 0 356574 800
rect 357346 0 357402 800
rect 358174 0 358230 800
rect 359002 0 359058 800
rect 359830 0 359886 800
rect 360658 0 360714 800
rect 361486 0 361542 800
rect 362314 0 362370 800
rect 363142 0 363198 800
rect 363970 0 364026 800
rect 364798 0 364854 800
rect 365626 0 365682 800
rect 366454 0 366510 800
rect 367282 0 367338 800
rect 368110 0 368166 800
rect 368938 0 368994 800
rect 369766 0 369822 800
rect 370594 0 370650 800
rect 371422 0 371478 800
rect 372250 0 372306 800
rect 373078 0 373134 800
rect 373906 0 373962 800
rect 374734 0 374790 800
rect 375562 0 375618 800
rect 376390 0 376446 800
rect 377218 0 377274 800
rect 378046 0 378102 800
rect 378874 0 378930 800
rect 379702 0 379758 800
rect 380530 0 380586 800
rect 381358 0 381414 800
rect 382186 0 382242 800
rect 383014 0 383070 800
rect 383842 0 383898 800
rect 384670 0 384726 800
rect 385498 0 385554 800
rect 386326 0 386382 800
rect 387154 0 387210 800
rect 387982 0 388038 800
rect 388810 0 388866 800
rect 389638 0 389694 800
rect 390466 0 390522 800
rect 391294 0 391350 800
rect 392122 0 392178 800
rect 392950 0 393006 800
rect 393778 0 393834 800
rect 394606 0 394662 800
rect 395434 0 395490 800
rect 396262 0 396318 800
rect 397090 0 397146 800
rect 397918 0 397974 800
rect 398746 0 398802 800
rect 399574 0 399630 800
rect 400402 0 400458 800
rect 401230 0 401286 800
rect 402058 0 402114 800
rect 402886 0 402942 800
rect 403714 0 403770 800
rect 404542 0 404598 800
rect 405370 0 405426 800
rect 406198 0 406254 800
rect 407026 0 407082 800
rect 407854 0 407910 800
rect 408682 0 408738 800
rect 409510 0 409566 800
rect 410338 0 410394 800
rect 411166 0 411222 800
rect 411994 0 412050 800
rect 412822 0 412878 800
rect 413650 0 413706 800
rect 414478 0 414534 800
rect 415306 0 415362 800
rect 416134 0 416190 800
rect 416962 0 417018 800
rect 417790 0 417846 800
rect 418618 0 418674 800
rect 419446 0 419502 800
rect 420274 0 420330 800
rect 421102 0 421158 800
rect 421930 0 421986 800
rect 422758 0 422814 800
rect 423586 0 423642 800
<< obsm2 >>
rect 938 856 438638 437413
rect 938 734 16154 856
rect 16322 734 16982 856
rect 17150 734 17810 856
rect 17978 734 18638 856
rect 18806 734 19466 856
rect 19634 734 20294 856
rect 20462 734 21122 856
rect 21290 734 21950 856
rect 22118 734 22778 856
rect 22946 734 23606 856
rect 23774 734 24434 856
rect 24602 734 25262 856
rect 25430 734 26090 856
rect 26258 734 26918 856
rect 27086 734 27746 856
rect 27914 734 28574 856
rect 28742 734 29402 856
rect 29570 734 30230 856
rect 30398 734 31058 856
rect 31226 734 31886 856
rect 32054 734 32714 856
rect 32882 734 33542 856
rect 33710 734 34370 856
rect 34538 734 35198 856
rect 35366 734 36026 856
rect 36194 734 36854 856
rect 37022 734 37682 856
rect 37850 734 38510 856
rect 38678 734 39338 856
rect 39506 734 40166 856
rect 40334 734 40994 856
rect 41162 734 41822 856
rect 41990 734 42650 856
rect 42818 734 43478 856
rect 43646 734 44306 856
rect 44474 734 45134 856
rect 45302 734 45962 856
rect 46130 734 46790 856
rect 46958 734 47618 856
rect 47786 734 48446 856
rect 48614 734 49274 856
rect 49442 734 50102 856
rect 50270 734 50930 856
rect 51098 734 51758 856
rect 51926 734 52586 856
rect 52754 734 53414 856
rect 53582 734 54242 856
rect 54410 734 55070 856
rect 55238 734 55898 856
rect 56066 734 56726 856
rect 56894 734 57554 856
rect 57722 734 58382 856
rect 58550 734 59210 856
rect 59378 734 60038 856
rect 60206 734 60866 856
rect 61034 734 61694 856
rect 61862 734 62522 856
rect 62690 734 63350 856
rect 63518 734 64178 856
rect 64346 734 65006 856
rect 65174 734 65834 856
rect 66002 734 66662 856
rect 66830 734 67490 856
rect 67658 734 68318 856
rect 68486 734 69146 856
rect 69314 734 69974 856
rect 70142 734 70802 856
rect 70970 734 71630 856
rect 71798 734 72458 856
rect 72626 734 73286 856
rect 73454 734 74114 856
rect 74282 734 74942 856
rect 75110 734 75770 856
rect 75938 734 76598 856
rect 76766 734 77426 856
rect 77594 734 78254 856
rect 78422 734 79082 856
rect 79250 734 79910 856
rect 80078 734 80738 856
rect 80906 734 81566 856
rect 81734 734 82394 856
rect 82562 734 83222 856
rect 83390 734 84050 856
rect 84218 734 84878 856
rect 85046 734 85706 856
rect 85874 734 86534 856
rect 86702 734 87362 856
rect 87530 734 88190 856
rect 88358 734 89018 856
rect 89186 734 89846 856
rect 90014 734 90674 856
rect 90842 734 91502 856
rect 91670 734 92330 856
rect 92498 734 93158 856
rect 93326 734 93986 856
rect 94154 734 94814 856
rect 94982 734 95642 856
rect 95810 734 96470 856
rect 96638 734 97298 856
rect 97466 734 98126 856
rect 98294 734 98954 856
rect 99122 734 99782 856
rect 99950 734 100610 856
rect 100778 734 101438 856
rect 101606 734 102266 856
rect 102434 734 103094 856
rect 103262 734 103922 856
rect 104090 734 104750 856
rect 104918 734 105578 856
rect 105746 734 106406 856
rect 106574 734 107234 856
rect 107402 734 108062 856
rect 108230 734 108890 856
rect 109058 734 109718 856
rect 109886 734 110546 856
rect 110714 734 111374 856
rect 111542 734 112202 856
rect 112370 734 113030 856
rect 113198 734 113858 856
rect 114026 734 114686 856
rect 114854 734 115514 856
rect 115682 734 116342 856
rect 116510 734 117170 856
rect 117338 734 117998 856
rect 118166 734 118826 856
rect 118994 734 119654 856
rect 119822 734 120482 856
rect 120650 734 121310 856
rect 121478 734 122138 856
rect 122306 734 122966 856
rect 123134 734 123794 856
rect 123962 734 124622 856
rect 124790 734 125450 856
rect 125618 734 126278 856
rect 126446 734 127106 856
rect 127274 734 127934 856
rect 128102 734 128762 856
rect 128930 734 129590 856
rect 129758 734 130418 856
rect 130586 734 131246 856
rect 131414 734 132074 856
rect 132242 734 132902 856
rect 133070 734 133730 856
rect 133898 734 134558 856
rect 134726 734 135386 856
rect 135554 734 136214 856
rect 136382 734 137042 856
rect 137210 734 137870 856
rect 138038 734 138698 856
rect 138866 734 139526 856
rect 139694 734 140354 856
rect 140522 734 141182 856
rect 141350 734 142010 856
rect 142178 734 142838 856
rect 143006 734 143666 856
rect 143834 734 144494 856
rect 144662 734 145322 856
rect 145490 734 146150 856
rect 146318 734 146978 856
rect 147146 734 147806 856
rect 147974 734 148634 856
rect 148802 734 149462 856
rect 149630 734 150290 856
rect 150458 734 151118 856
rect 151286 734 151946 856
rect 152114 734 152774 856
rect 152942 734 153602 856
rect 153770 734 154430 856
rect 154598 734 155258 856
rect 155426 734 156086 856
rect 156254 734 156914 856
rect 157082 734 157742 856
rect 157910 734 158570 856
rect 158738 734 159398 856
rect 159566 734 160226 856
rect 160394 734 161054 856
rect 161222 734 161882 856
rect 162050 734 162710 856
rect 162878 734 163538 856
rect 163706 734 164366 856
rect 164534 734 165194 856
rect 165362 734 166022 856
rect 166190 734 166850 856
rect 167018 734 167678 856
rect 167846 734 168506 856
rect 168674 734 169334 856
rect 169502 734 170162 856
rect 170330 734 170990 856
rect 171158 734 171818 856
rect 171986 734 172646 856
rect 172814 734 173474 856
rect 173642 734 174302 856
rect 174470 734 175130 856
rect 175298 734 175958 856
rect 176126 734 176786 856
rect 176954 734 177614 856
rect 177782 734 178442 856
rect 178610 734 179270 856
rect 179438 734 180098 856
rect 180266 734 180926 856
rect 181094 734 181754 856
rect 181922 734 182582 856
rect 182750 734 183410 856
rect 183578 734 184238 856
rect 184406 734 185066 856
rect 185234 734 185894 856
rect 186062 734 186722 856
rect 186890 734 187550 856
rect 187718 734 188378 856
rect 188546 734 189206 856
rect 189374 734 190034 856
rect 190202 734 190862 856
rect 191030 734 191690 856
rect 191858 734 192518 856
rect 192686 734 193346 856
rect 193514 734 194174 856
rect 194342 734 195002 856
rect 195170 734 195830 856
rect 195998 734 196658 856
rect 196826 734 197486 856
rect 197654 734 198314 856
rect 198482 734 199142 856
rect 199310 734 199970 856
rect 200138 734 200798 856
rect 200966 734 201626 856
rect 201794 734 202454 856
rect 202622 734 203282 856
rect 203450 734 204110 856
rect 204278 734 204938 856
rect 205106 734 205766 856
rect 205934 734 206594 856
rect 206762 734 207422 856
rect 207590 734 208250 856
rect 208418 734 209078 856
rect 209246 734 209906 856
rect 210074 734 210734 856
rect 210902 734 211562 856
rect 211730 734 212390 856
rect 212558 734 213218 856
rect 213386 734 214046 856
rect 214214 734 214874 856
rect 215042 734 215702 856
rect 215870 734 216530 856
rect 216698 734 217358 856
rect 217526 734 218186 856
rect 218354 734 219014 856
rect 219182 734 219842 856
rect 220010 734 220670 856
rect 220838 734 221498 856
rect 221666 734 222326 856
rect 222494 734 223154 856
rect 223322 734 223982 856
rect 224150 734 224810 856
rect 224978 734 225638 856
rect 225806 734 226466 856
rect 226634 734 227294 856
rect 227462 734 228122 856
rect 228290 734 228950 856
rect 229118 734 229778 856
rect 229946 734 230606 856
rect 230774 734 231434 856
rect 231602 734 232262 856
rect 232430 734 233090 856
rect 233258 734 233918 856
rect 234086 734 234746 856
rect 234914 734 235574 856
rect 235742 734 236402 856
rect 236570 734 237230 856
rect 237398 734 238058 856
rect 238226 734 238886 856
rect 239054 734 239714 856
rect 239882 734 240542 856
rect 240710 734 241370 856
rect 241538 734 242198 856
rect 242366 734 243026 856
rect 243194 734 243854 856
rect 244022 734 244682 856
rect 244850 734 245510 856
rect 245678 734 246338 856
rect 246506 734 247166 856
rect 247334 734 247994 856
rect 248162 734 248822 856
rect 248990 734 249650 856
rect 249818 734 250478 856
rect 250646 734 251306 856
rect 251474 734 252134 856
rect 252302 734 252962 856
rect 253130 734 253790 856
rect 253958 734 254618 856
rect 254786 734 255446 856
rect 255614 734 256274 856
rect 256442 734 257102 856
rect 257270 734 257930 856
rect 258098 734 258758 856
rect 258926 734 259586 856
rect 259754 734 260414 856
rect 260582 734 261242 856
rect 261410 734 262070 856
rect 262238 734 262898 856
rect 263066 734 263726 856
rect 263894 734 264554 856
rect 264722 734 265382 856
rect 265550 734 266210 856
rect 266378 734 267038 856
rect 267206 734 267866 856
rect 268034 734 268694 856
rect 268862 734 269522 856
rect 269690 734 270350 856
rect 270518 734 271178 856
rect 271346 734 272006 856
rect 272174 734 272834 856
rect 273002 734 273662 856
rect 273830 734 274490 856
rect 274658 734 275318 856
rect 275486 734 276146 856
rect 276314 734 276974 856
rect 277142 734 277802 856
rect 277970 734 278630 856
rect 278798 734 279458 856
rect 279626 734 280286 856
rect 280454 734 281114 856
rect 281282 734 281942 856
rect 282110 734 282770 856
rect 282938 734 283598 856
rect 283766 734 284426 856
rect 284594 734 285254 856
rect 285422 734 286082 856
rect 286250 734 286910 856
rect 287078 734 287738 856
rect 287906 734 288566 856
rect 288734 734 289394 856
rect 289562 734 290222 856
rect 290390 734 291050 856
rect 291218 734 291878 856
rect 292046 734 292706 856
rect 292874 734 293534 856
rect 293702 734 294362 856
rect 294530 734 295190 856
rect 295358 734 296018 856
rect 296186 734 296846 856
rect 297014 734 297674 856
rect 297842 734 298502 856
rect 298670 734 299330 856
rect 299498 734 300158 856
rect 300326 734 300986 856
rect 301154 734 301814 856
rect 301982 734 302642 856
rect 302810 734 303470 856
rect 303638 734 304298 856
rect 304466 734 305126 856
rect 305294 734 305954 856
rect 306122 734 306782 856
rect 306950 734 307610 856
rect 307778 734 308438 856
rect 308606 734 309266 856
rect 309434 734 310094 856
rect 310262 734 310922 856
rect 311090 734 311750 856
rect 311918 734 312578 856
rect 312746 734 313406 856
rect 313574 734 314234 856
rect 314402 734 315062 856
rect 315230 734 315890 856
rect 316058 734 316718 856
rect 316886 734 317546 856
rect 317714 734 318374 856
rect 318542 734 319202 856
rect 319370 734 320030 856
rect 320198 734 320858 856
rect 321026 734 321686 856
rect 321854 734 322514 856
rect 322682 734 323342 856
rect 323510 734 324170 856
rect 324338 734 324998 856
rect 325166 734 325826 856
rect 325994 734 326654 856
rect 326822 734 327482 856
rect 327650 734 328310 856
rect 328478 734 329138 856
rect 329306 734 329966 856
rect 330134 734 330794 856
rect 330962 734 331622 856
rect 331790 734 332450 856
rect 332618 734 333278 856
rect 333446 734 334106 856
rect 334274 734 334934 856
rect 335102 734 335762 856
rect 335930 734 336590 856
rect 336758 734 337418 856
rect 337586 734 338246 856
rect 338414 734 339074 856
rect 339242 734 339902 856
rect 340070 734 340730 856
rect 340898 734 341558 856
rect 341726 734 342386 856
rect 342554 734 343214 856
rect 343382 734 344042 856
rect 344210 734 344870 856
rect 345038 734 345698 856
rect 345866 734 346526 856
rect 346694 734 347354 856
rect 347522 734 348182 856
rect 348350 734 349010 856
rect 349178 734 349838 856
rect 350006 734 350666 856
rect 350834 734 351494 856
rect 351662 734 352322 856
rect 352490 734 353150 856
rect 353318 734 353978 856
rect 354146 734 354806 856
rect 354974 734 355634 856
rect 355802 734 356462 856
rect 356630 734 357290 856
rect 357458 734 358118 856
rect 358286 734 358946 856
rect 359114 734 359774 856
rect 359942 734 360602 856
rect 360770 734 361430 856
rect 361598 734 362258 856
rect 362426 734 363086 856
rect 363254 734 363914 856
rect 364082 734 364742 856
rect 364910 734 365570 856
rect 365738 734 366398 856
rect 366566 734 367226 856
rect 367394 734 368054 856
rect 368222 734 368882 856
rect 369050 734 369710 856
rect 369878 734 370538 856
rect 370706 734 371366 856
rect 371534 734 372194 856
rect 372362 734 373022 856
rect 373190 734 373850 856
rect 374018 734 374678 856
rect 374846 734 375506 856
rect 375674 734 376334 856
rect 376502 734 377162 856
rect 377330 734 377990 856
rect 378158 734 378818 856
rect 378986 734 379646 856
rect 379814 734 380474 856
rect 380642 734 381302 856
rect 381470 734 382130 856
rect 382298 734 382958 856
rect 383126 734 383786 856
rect 383954 734 384614 856
rect 384782 734 385442 856
rect 385610 734 386270 856
rect 386438 734 387098 856
rect 387266 734 387926 856
rect 388094 734 388754 856
rect 388922 734 389582 856
rect 389750 734 390410 856
rect 390578 734 391238 856
rect 391406 734 392066 856
rect 392234 734 392894 856
rect 393062 734 393722 856
rect 393890 734 394550 856
rect 394718 734 395378 856
rect 395546 734 396206 856
rect 396374 734 397034 856
rect 397202 734 397862 856
rect 398030 734 398690 856
rect 398858 734 399518 856
rect 399686 734 400346 856
rect 400514 734 401174 856
rect 401342 734 402002 856
rect 402170 734 402830 856
rect 402998 734 403658 856
rect 403826 734 404486 856
rect 404654 734 405314 856
rect 405482 734 406142 856
rect 406310 734 406970 856
rect 407138 734 407798 856
rect 407966 734 408626 856
rect 408794 734 409454 856
rect 409622 734 410282 856
rect 410450 734 411110 856
rect 411278 734 411938 856
rect 412106 734 412766 856
rect 412934 734 413594 856
rect 413762 734 414422 856
rect 414590 734 415250 856
rect 415418 734 416078 856
rect 416246 734 416906 856
rect 417074 734 417734 856
rect 417902 734 418562 856
rect 418730 734 419390 856
rect 419558 734 420218 856
rect 420386 734 421046 856
rect 421214 734 421874 856
rect 422042 734 422702 856
rect 422870 734 423530 856
rect 423698 734 438638 856
<< metal3 >>
rect 0 433032 800 433152
rect 439200 433032 440000 433152
rect 0 425416 800 425536
rect 439200 425416 440000 425536
rect 0 417800 800 417920
rect 439200 417800 440000 417920
rect 0 410184 800 410304
rect 439200 410184 440000 410304
rect 0 402568 800 402688
rect 439200 402568 440000 402688
rect 0 394952 800 395072
rect 439200 394952 440000 395072
rect 0 387336 800 387456
rect 439200 387336 440000 387456
rect 0 379720 800 379840
rect 439200 379720 440000 379840
rect 0 372104 800 372224
rect 439200 372104 440000 372224
rect 0 364488 800 364608
rect 439200 364488 440000 364608
rect 0 356872 800 356992
rect 439200 356872 440000 356992
rect 0 349256 800 349376
rect 439200 349256 440000 349376
rect 0 341640 800 341760
rect 439200 341640 440000 341760
rect 0 334024 800 334144
rect 439200 334024 440000 334144
rect 0 326408 800 326528
rect 439200 326408 440000 326528
rect 0 318792 800 318912
rect 439200 318792 440000 318912
rect 0 311176 800 311296
rect 439200 311176 440000 311296
rect 0 303560 800 303680
rect 439200 303560 440000 303680
rect 0 295944 800 296064
rect 439200 295944 440000 296064
rect 0 288328 800 288448
rect 439200 288328 440000 288448
rect 0 280712 800 280832
rect 439200 280712 440000 280832
rect 0 273096 800 273216
rect 439200 273096 440000 273216
rect 0 265480 800 265600
rect 439200 265480 440000 265600
rect 0 257864 800 257984
rect 439200 257864 440000 257984
rect 0 250248 800 250368
rect 439200 250248 440000 250368
rect 0 242632 800 242752
rect 439200 242632 440000 242752
rect 0 235016 800 235136
rect 439200 235016 440000 235136
rect 0 227400 800 227520
rect 439200 227400 440000 227520
rect 0 219784 800 219904
rect 439200 219784 440000 219904
rect 0 212168 800 212288
rect 439200 212168 440000 212288
rect 0 204552 800 204672
rect 439200 204552 440000 204672
rect 0 196936 800 197056
rect 439200 196936 440000 197056
rect 0 189320 800 189440
rect 439200 189320 440000 189440
rect 0 181704 800 181824
rect 439200 181704 440000 181824
rect 0 174088 800 174208
rect 439200 174088 440000 174208
rect 0 166472 800 166592
rect 439200 166472 440000 166592
rect 0 158856 800 158976
rect 439200 158856 440000 158976
rect 0 151240 800 151360
rect 439200 151240 440000 151360
rect 0 143624 800 143744
rect 439200 143624 440000 143744
rect 0 136008 800 136128
rect 439200 136008 440000 136128
rect 0 128392 800 128512
rect 439200 128392 440000 128512
rect 0 120776 800 120896
rect 439200 120776 440000 120896
rect 0 113160 800 113280
rect 439200 113160 440000 113280
rect 0 105544 800 105664
rect 439200 105544 440000 105664
rect 0 97928 800 98048
rect 439200 97928 440000 98048
rect 0 90312 800 90432
rect 439200 90312 440000 90432
rect 0 82696 800 82816
rect 439200 82696 440000 82816
rect 0 75080 800 75200
rect 439200 75080 440000 75200
rect 0 67464 800 67584
rect 439200 67464 440000 67584
rect 0 59848 800 59968
rect 439200 59848 440000 59968
rect 0 52232 800 52352
rect 439200 52232 440000 52352
rect 0 44616 800 44736
rect 439200 44616 440000 44736
rect 0 37000 800 37120
rect 439200 37000 440000 37120
rect 0 29384 800 29504
rect 439200 29384 440000 29504
rect 0 21768 800 21888
rect 439200 21768 440000 21888
rect 0 14152 800 14272
rect 439200 14152 440000 14272
rect 0 6536 800 6656
rect 439200 6536 440000 6656
<< obsm3 >>
rect 798 433232 439200 437409
rect 880 432952 439120 433232
rect 798 425616 439200 432952
rect 880 425336 439120 425616
rect 798 418000 439200 425336
rect 880 417720 439120 418000
rect 798 410384 439200 417720
rect 880 410104 439120 410384
rect 798 402768 439200 410104
rect 880 402488 439120 402768
rect 798 395152 439200 402488
rect 880 394872 439120 395152
rect 798 387536 439200 394872
rect 880 387256 439120 387536
rect 798 379920 439200 387256
rect 880 379640 439120 379920
rect 798 372304 439200 379640
rect 880 372024 439120 372304
rect 798 364688 439200 372024
rect 880 364408 439120 364688
rect 798 357072 439200 364408
rect 880 356792 439120 357072
rect 798 349456 439200 356792
rect 880 349176 439120 349456
rect 798 341840 439200 349176
rect 880 341560 439120 341840
rect 798 334224 439200 341560
rect 880 333944 439120 334224
rect 798 326608 439200 333944
rect 880 326328 439120 326608
rect 798 318992 439200 326328
rect 880 318712 439120 318992
rect 798 311376 439200 318712
rect 880 311096 439120 311376
rect 798 303760 439200 311096
rect 880 303480 439120 303760
rect 798 296144 439200 303480
rect 880 295864 439120 296144
rect 798 288528 439200 295864
rect 880 288248 439120 288528
rect 798 280912 439200 288248
rect 880 280632 439120 280912
rect 798 273296 439200 280632
rect 880 273016 439120 273296
rect 798 265680 439200 273016
rect 880 265400 439120 265680
rect 798 258064 439200 265400
rect 880 257784 439120 258064
rect 798 250448 439200 257784
rect 880 250168 439120 250448
rect 798 242832 439200 250168
rect 880 242552 439120 242832
rect 798 235216 439200 242552
rect 880 234936 439120 235216
rect 798 227600 439200 234936
rect 880 227320 439120 227600
rect 798 219984 439200 227320
rect 880 219704 439120 219984
rect 798 212368 439200 219704
rect 880 212088 439120 212368
rect 798 204752 439200 212088
rect 880 204472 439120 204752
rect 798 197136 439200 204472
rect 880 196856 439120 197136
rect 798 189520 439200 196856
rect 880 189240 439120 189520
rect 798 181904 439200 189240
rect 880 181624 439120 181904
rect 798 174288 439200 181624
rect 880 174008 439120 174288
rect 798 166672 439200 174008
rect 880 166392 439120 166672
rect 798 159056 439200 166392
rect 880 158776 439120 159056
rect 798 151440 439200 158776
rect 880 151160 439120 151440
rect 798 143824 439200 151160
rect 880 143544 439120 143824
rect 798 136208 439200 143544
rect 880 135928 439120 136208
rect 798 128592 439200 135928
rect 880 128312 439120 128592
rect 798 120976 439200 128312
rect 880 120696 439120 120976
rect 798 113360 439200 120696
rect 880 113080 439120 113360
rect 798 105744 439200 113080
rect 880 105464 439120 105744
rect 798 98128 439200 105464
rect 880 97848 439120 98128
rect 798 90512 439200 97848
rect 880 90232 439120 90512
rect 798 82896 439200 90232
rect 880 82616 439120 82896
rect 798 75280 439200 82616
rect 880 75000 439120 75280
rect 798 67664 439200 75000
rect 880 67384 439120 67664
rect 798 60048 439200 67384
rect 880 59768 439120 60048
rect 798 52432 439200 59768
rect 880 52152 439120 52432
rect 798 44816 439200 52152
rect 880 44536 439120 44816
rect 798 37200 439200 44536
rect 880 36920 439120 37200
rect 798 29584 439200 36920
rect 880 29304 439120 29584
rect 798 21968 439200 29304
rect 880 21688 439120 21968
rect 798 14352 439200 21688
rect 880 14072 439120 14352
rect 798 6736 439200 14072
rect 880 6456 439120 6736
rect 798 1939 439200 6456
<< metal4 >>
rect 4208 2128 4528 437424
rect 19568 2128 19888 437424
rect 34928 2128 35248 437424
rect 50288 2128 50608 437424
rect 65648 2128 65968 437424
rect 81008 2128 81328 437424
rect 96368 2128 96688 437424
rect 111728 2128 112048 437424
rect 127088 2128 127408 437424
rect 142448 2128 142768 437424
rect 157808 2128 158128 437424
rect 173168 2128 173488 437424
rect 188528 2128 188848 437424
rect 203888 2128 204208 437424
rect 219248 2128 219568 437424
rect 234608 2128 234928 437424
rect 249968 2128 250288 437424
rect 265328 2128 265648 437424
rect 280688 2128 281008 437424
rect 296048 2128 296368 437424
rect 311408 2128 311728 437424
rect 326768 2128 327088 437424
rect 342128 2128 342448 437424
rect 357488 2128 357808 437424
rect 372848 2128 373168 437424
rect 388208 2128 388528 437424
rect 403568 2128 403888 437424
rect 418928 2128 419248 437424
rect 434288 2128 434608 437424
<< obsm4 >>
rect 88747 6699 96288 329901
rect 96768 6699 111648 329901
rect 112128 6699 127008 329901
rect 127488 6699 142368 329901
rect 142848 6699 157728 329901
rect 158208 6699 173088 329901
rect 173568 6699 188448 329901
rect 188928 6699 203808 329901
rect 204288 6699 219168 329901
rect 219648 6699 234528 329901
rect 235008 6699 249888 329901
rect 250368 6699 265248 329901
rect 265728 6699 280608 329901
rect 281088 6699 295968 329901
rect 296448 6699 311328 329901
rect 311808 6699 314949 329901
<< labels >>
rlabel metal3 s 439200 6536 440000 6656 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 439200 235016 440000 235136 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 439200 257864 440000 257984 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 439200 280712 440000 280832 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 439200 303560 440000 303680 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 439200 326408 440000 326528 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 439200 349256 440000 349376 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 439200 372104 440000 372224 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 439200 394952 440000 395072 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 439200 417800 440000 417920 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 433032 800 433152 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 439200 29384 440000 29504 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 410184 800 410304 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 387336 800 387456 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 0 364488 800 364608 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 0 341640 800 341760 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 318792 800 318912 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 295944 800 296064 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 273096 800 273216 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 250248 800 250368 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 227400 800 227520 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 204552 800 204672 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 439200 52232 440000 52352 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 181704 800 181824 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 158856 800 158976 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 439200 75080 440000 75200 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 439200 97928 440000 98048 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 439200 120776 440000 120896 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 439200 143624 440000 143744 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 439200 166472 440000 166592 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 439200 189320 440000 189440 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 439200 212168 440000 212288 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 439200 21768 440000 21888 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 439200 250248 440000 250368 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 439200 273096 440000 273216 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 439200 295944 440000 296064 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 439200 318792 440000 318912 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 439200 341640 440000 341760 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 439200 364488 440000 364608 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 439200 387336 440000 387456 6 io_oeb[16]
port 46 nsew signal output
rlabel metal3 s 439200 410184 440000 410304 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 439200 433032 440000 433152 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 417800 800 417920 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 439200 44616 440000 44736 6 io_oeb[1]
port 50 nsew signal output
rlabel metal3 s 0 394952 800 395072 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 0 372104 800 372224 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 0 349256 800 349376 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 326408 800 326528 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 303560 800 303680 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 280712 800 280832 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 257864 800 257984 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 235016 800 235136 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 212168 800 212288 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 189320 800 189440 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 439200 67464 440000 67584 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 166472 800 166592 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 143624 800 143744 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 120776 800 120896 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 75080 800 75200 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 439200 90312 440000 90432 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 439200 113160 440000 113280 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 439200 136008 440000 136128 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 439200 158856 440000 158976 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 439200 181704 440000 181824 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 439200 204552 440000 204672 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 439200 227400 440000 227520 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 439200 14152 440000 14272 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 439200 242632 440000 242752 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 439200 265480 440000 265600 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 439200 288328 440000 288448 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 439200 311176 440000 311296 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 439200 334024 440000 334144 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 439200 356872 440000 356992 6 io_out[15]
port 83 nsew signal output
rlabel metal3 s 439200 379720 440000 379840 6 io_out[16]
port 84 nsew signal output
rlabel metal3 s 439200 402568 440000 402688 6 io_out[17]
port 85 nsew signal output
rlabel metal3 s 439200 425416 440000 425536 6 io_out[18]
port 86 nsew signal output
rlabel metal3 s 0 425416 800 425536 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 439200 37000 440000 37120 6 io_out[1]
port 88 nsew signal output
rlabel metal3 s 0 402568 800 402688 6 io_out[20]
port 89 nsew signal output
rlabel metal3 s 0 379720 800 379840 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 0 356872 800 356992 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 0 334024 800 334144 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 311176 800 311296 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 288328 800 288448 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 265480 800 265600 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 242632 800 242752 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 219784 800 219904 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 196936 800 197056 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 439200 59848 440000 59968 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 151240 800 151360 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 439200 82696 440000 82816 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 439200 105544 440000 105664 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 439200 128392 440000 128512 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 439200 151240 440000 151360 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 439200 174088 440000 174208 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 439200 196936 440000 197056 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 439200 219784 440000 219904 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 421930 0 421986 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 422758 0 422814 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 423586 0 423642 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 352378 0 352434 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 354862 0 354918 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 357346 0 357402 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 359830 0 359886 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 362314 0 362370 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 364798 0 364854 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 367282 0 367338 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 369766 0 369822 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 372250 0 372306 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 374734 0 374790 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 377218 0 377274 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 379702 0 379758 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 382186 0 382242 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 384670 0 384726 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 387154 0 387210 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 389638 0 389694 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 392122 0 392178 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 394606 0 394662 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 397090 0 397146 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 402058 0 402114 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 404542 0 404598 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 407026 0 407082 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 409510 0 409566 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 411994 0 412050 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 414478 0 414534 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 416962 0 417018 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 419446 0 419502 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 158626 0 158682 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 166078 0 166134 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 176014 0 176070 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 190918 0 190974 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 193402 0 193458 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 200854 0 200910 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 205822 0 205878 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 210790 0 210846 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 238114 0 238170 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 240598 0 240654 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 243082 0 243138 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 250534 0 250590 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 253018 0 253074 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 255502 0 255558 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 260470 0 260526 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 265438 0 265494 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 267922 0 267978 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 270406 0 270462 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 280342 0 280398 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 285310 0 285366 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 287794 0 287850 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 290278 0 290334 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 292762 0 292818 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 295246 0 295302 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 297730 0 297786 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 300214 0 300270 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 302698 0 302754 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 305182 0 305238 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 310150 0 310206 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 312634 0 312690 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 320086 0 320142 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 322570 0 322626 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 327538 0 327594 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 330022 0 330078 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 332506 0 332562 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 334990 0 335046 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 337474 0 337530 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 339958 0 340014 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 342442 0 342498 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 344926 0 344982 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 347410 0 347466 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 349894 0 349950 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 355690 0 355746 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 358174 0 358230 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 360658 0 360714 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 363142 0 363198 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 365626 0 365682 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 368110 0 368166 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 370594 0 370650 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 373078 0 373134 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 375562 0 375618 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 129646 0 129702 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 378046 0 378102 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 380530 0 380586 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 383014 0 383070 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 385498 0 385554 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 387982 0 388038 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 390466 0 390522 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 392950 0 393006 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 395434 0 395490 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 397918 0 397974 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 400402 0 400458 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 402886 0 402942 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 405370 0 405426 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 410338 0 410394 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 412822 0 412878 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 415306 0 415362 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 417790 0 417846 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 420274 0 420330 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 142066 0 142122 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 107290 0 107346 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 154486 0 154542 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 159454 0 159510 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 166906 0 166962 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 169390 0 169446 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 171874 0 171930 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 181810 0 181866 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 184294 0 184350 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 189262 0 189318 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 209134 0 209190 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 211618 0 211674 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 226522 0 226578 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 229006 0 229062 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 233974 0 234030 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 238942 0 238998 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 241426 0 241482 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 243910 0 243966 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 246394 0 246450 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 251362 0 251418 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 253846 0 253902 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 256330 0 256386 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 258814 0 258870 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 261298 0 261354 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 268750 0 268806 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 271234 0 271290 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 273718 0 273774 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 276202 0 276258 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 278686 0 278742 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 281170 0 281226 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 286138 0 286194 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 288622 0 288678 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 291106 0 291162 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 293590 0 293646 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 296074 0 296130 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 122194 0 122250 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 303526 0 303582 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 306010 0 306066 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 308494 0 308550 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 310978 0 311034 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 313462 0 313518 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 320914 0 320970 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 323398 0 323454 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 325882 0 325938 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 330850 0 330906 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 335818 0 335874 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 338302 0 338358 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 340786 0 340842 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 343270 0 343326 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 345754 0 345810 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 348238 0 348294 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 350722 0 350778 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 356518 0 356574 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 361486 0 361542 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 363970 0 364026 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 366454 0 366510 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 368938 0 368994 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 371422 0 371478 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 373906 0 373962 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 376390 0 376446 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 378874 0 378930 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 381358 0 381414 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 383842 0 383898 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 386326 0 386382 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 388810 0 388866 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 391294 0 391350 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 393778 0 393834 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 396262 0 396318 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 398746 0 398802 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 401230 0 401286 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 403714 0 403770 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 406198 0 406254 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 408682 0 408738 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 413650 0 413706 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 416134 0 416190 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 418618 0 418674 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 421102 0 421158 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 147862 0 147918 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 155314 0 155370 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 180154 0 180210 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 200026 0 200082 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 209962 0 210018 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 222382 0 222438 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 224866 0 224922 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 227350 0 227406 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 229834 0 229890 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 244738 0 244794 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 249706 0 249762 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 254674 0 254730 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 257158 0 257214 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 267094 0 267150 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 269578 0 269634 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 272062 0 272118 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 277030 0 277086 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 279514 0 279570 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 281998 0 282054 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 289450 0 289506 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 291934 0 291990 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 294418 0 294474 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 296902 0 296958 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 301870 0 301926 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 304354 0 304410 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 306838 0 306894 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 309322 0 309378 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 314290 0 314346 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 321742 0 321798 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 326710 0 326766 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 329194 0 329250 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 331678 0 331734 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 334162 0 334218 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 336646 0 336702 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 339130 0 339186 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 341614 0 341670 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 344098 0 344154 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 346582 0 346638 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 349066 0 349122 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 351550 0 351606 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 437424 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 437424 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 16210 0 16266 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 71686 0 71742 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 440000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 137760592
string GDS_FILE /ux1/users/asinghan/caravel_user_project-mpw-9i/openlane/user_proj_example/runs/24_05_29_02_05/results/signoff/user_proj_example.magic.gds
string GDS_START 1875756
<< end >>

