magic
tech sky130A
magscale 1 2
timestamp 1682005840
<< viali >>
rect 949 4097 983 4131
rect 1593 4097 1627 4131
rect 1501 3485 1535 3519
rect 2513 3485 2547 3519
rect 1225 3009 1259 3043
rect 1685 3009 1719 3043
rect 1041 2397 1075 2431
rect 1041 1921 1075 1955
rect 1777 1921 1811 1955
rect 2421 1921 2455 1955
rect 949 1309 983 1343
rect 1593 1309 1627 1343
rect 2329 1309 2363 1343
<< metal1 >>
rect 460 4378 3220 4400
rect 460 4326 2698 4378
rect 2750 4326 2762 4378
rect 2814 4326 2826 4378
rect 2878 4326 2890 4378
rect 2942 4326 3220 4378
rect 460 4304 3220 4326
rect 937 4128 995 4137
rect 1121 4128 1179 4137
rect 1581 4128 1639 4137
rect 1765 4128 1823 4137
rect 937 4100 1179 4128
rect 937 4091 995 4100
rect 1121 4091 1179 4100
rect 1373 4100 1823 4128
rect 1136 4004 1164 4091
rect 1118 3952 1124 4004
rect 1176 3952 1182 4004
rect 1210 3884 1216 3936
rect 1268 3924 1274 3936
rect 1373 3924 1401 4100
rect 1581 4091 1639 4100
rect 1765 4091 1823 4100
rect 1268 3896 1401 3924
rect 1268 3884 1274 3896
rect 460 3834 3220 3856
rect 460 3782 818 3834
rect 870 3782 882 3834
rect 934 3782 946 3834
rect 998 3782 1010 3834
rect 1062 3782 3220 3834
rect 460 3760 3220 3782
rect 1394 3680 1400 3732
rect 1452 3680 1458 3732
rect 1415 3516 1443 3680
rect 1486 3612 1492 3664
rect 1544 3652 1550 3664
rect 1544 3624 2112 3652
rect 1544 3612 1550 3624
rect 1489 3516 1547 3525
rect 1673 3516 1731 3525
rect 1415 3488 1731 3516
rect 2084 3516 2112 3624
rect 2317 3516 2375 3525
rect 2501 3516 2559 3525
rect 2084 3488 2559 3516
rect 1489 3479 1547 3488
rect 1673 3479 1731 3488
rect 2317 3479 2375 3488
rect 2501 3479 2559 3488
rect 460 3290 3220 3312
rect 460 3238 2698 3290
rect 2750 3238 2762 3290
rect 2814 3238 2826 3290
rect 2878 3238 2890 3290
rect 2942 3238 3220 3290
rect 460 3216 3220 3238
rect 658 3136 664 3188
rect 716 3176 722 3188
rect 716 3148 894 3176
rect 716 3136 722 3148
rect 866 3040 894 3148
rect 1029 3040 1087 3049
rect 1213 3040 1271 3049
rect 1673 3040 1731 3049
rect 1857 3040 1915 3049
rect 866 3012 1271 3040
rect 1029 3003 1087 3012
rect 1213 3003 1271 3012
rect 1403 3012 1915 3040
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 1403 2904 1431 3012
rect 1673 3003 1731 3012
rect 1857 3003 1915 3012
rect 1176 2876 1431 2904
rect 1176 2864 1182 2876
rect 460 2746 3220 2768
rect 460 2694 818 2746
rect 870 2694 882 2746
rect 934 2694 946 2746
rect 998 2694 1010 2746
rect 1062 2694 3220 2746
rect 460 2672 3220 2694
rect 1118 2592 1124 2644
rect 1176 2592 1182 2644
rect 1029 2428 1087 2437
rect 1133 2428 1161 2592
rect 1213 2428 1271 2437
rect 1029 2400 1271 2428
rect 1029 2391 1087 2400
rect 1213 2391 1271 2400
rect 460 2202 3220 2224
rect 460 2150 2698 2202
rect 2750 2150 2762 2202
rect 2814 2150 2826 2202
rect 2878 2150 2890 2202
rect 2942 2150 3220 2202
rect 460 2128 3220 2150
rect 1029 1952 1087 1961
rect 1118 1952 1124 1964
rect 1029 1924 1124 1952
rect 1029 1915 1087 1924
rect 1118 1912 1124 1924
rect 1176 1952 1182 1964
rect 1213 1952 1271 1961
rect 1176 1924 1271 1952
rect 1176 1912 1182 1924
rect 1213 1915 1271 1924
rect 1302 1912 1308 1964
rect 1360 1952 1366 1964
rect 1765 1952 1823 1961
rect 1949 1952 2007 1961
rect 2409 1952 2467 1961
rect 2593 1952 2651 1961
rect 1360 1924 2007 1952
rect 1360 1912 1366 1924
rect 1765 1915 1823 1924
rect 1949 1915 2007 1924
rect 2244 1924 2651 1952
rect 566 1776 572 1828
rect 624 1816 630 1828
rect 2244 1816 2272 1924
rect 2409 1915 2467 1924
rect 2593 1915 2651 1924
rect 624 1788 2272 1816
rect 624 1776 630 1788
rect 460 1658 3220 1680
rect 460 1606 818 1658
rect 870 1606 882 1658
rect 934 1606 946 1658
rect 998 1606 1010 1658
rect 1062 1606 3220 1658
rect 460 1584 3220 1606
rect 1210 1504 1216 1556
rect 1268 1544 1274 1556
rect 1268 1516 2012 1544
rect 1268 1504 1274 1516
rect 1118 1436 1124 1488
rect 1176 1476 1182 1488
rect 1176 1448 1475 1476
rect 1176 1436 1182 1448
rect 658 1368 664 1420
rect 716 1408 722 1420
rect 716 1380 855 1408
rect 716 1368 722 1380
rect 827 1340 855 1380
rect 937 1340 995 1349
rect 1121 1340 1179 1349
rect 827 1312 1179 1340
rect 1447 1340 1475 1448
rect 1581 1340 1639 1349
rect 1765 1340 1823 1349
rect 1447 1312 1823 1340
rect 1984 1340 2012 1516
rect 2317 1340 2375 1349
rect 2501 1340 2559 1349
rect 1984 1312 2559 1340
rect 937 1303 995 1312
rect 1121 1303 1179 1312
rect 1581 1303 1639 1312
rect 1765 1303 1823 1312
rect 2317 1303 2375 1312
rect 2501 1303 2559 1312
rect 460 1114 3220 1136
rect 460 1062 2698 1114
rect 2750 1062 2762 1114
rect 2814 1062 2826 1114
rect 2878 1062 2890 1114
rect 2942 1062 3220 1114
rect 460 1040 3220 1062
<< via1 >>
rect 2698 4326 2750 4378
rect 2762 4326 2814 4378
rect 2826 4326 2878 4378
rect 2890 4326 2942 4378
rect 1124 3952 1176 4004
rect 1216 3884 1268 3936
rect 818 3782 870 3834
rect 882 3782 934 3834
rect 946 3782 998 3834
rect 1010 3782 1062 3834
rect 1400 3680 1452 3732
rect 1492 3612 1544 3664
rect 2698 3238 2750 3290
rect 2762 3238 2814 3290
rect 2826 3238 2878 3290
rect 2890 3238 2942 3290
rect 664 3136 716 3188
rect 1124 2864 1176 2916
rect 818 2694 870 2746
rect 882 2694 934 2746
rect 946 2694 998 2746
rect 1010 2694 1062 2746
rect 1124 2592 1176 2644
rect 2698 2150 2750 2202
rect 2762 2150 2814 2202
rect 2826 2150 2878 2202
rect 2890 2150 2942 2202
rect 1124 1912 1176 1964
rect 1308 1912 1360 1964
rect 572 1776 624 1828
rect 818 1606 870 1658
rect 882 1606 934 1658
rect 946 1606 998 1658
rect 1010 1606 1062 1658
rect 1216 1504 1268 1556
rect 1124 1436 1176 1488
rect 664 1368 716 1420
rect 2698 1062 2750 1114
rect 2762 1062 2814 1114
rect 2826 1062 2878 1114
rect 2890 1062 2942 1114
<< metal2 >>
rect 754 5114 810 6200
rect 1122 5114 1178 6200
rect 754 5086 1072 5114
rect 754 5000 810 5086
rect 1044 4570 1072 5086
rect 1122 5086 1348 5114
rect 1122 5000 1178 5086
rect 1320 4706 1348 5086
rect 1320 4678 1440 4706
rect 1044 4542 1348 4570
rect 662 4448 718 4457
rect 662 4383 718 4392
rect 676 3194 704 4383
rect 800 3834 1080 4400
rect 1122 4040 1178 4049
rect 1122 3975 1124 3984
rect 1176 3975 1178 3984
rect 1124 3946 1176 3952
rect 1216 3936 1268 3942
rect 1216 3878 1268 3884
rect 800 3782 818 3834
rect 870 3782 882 3834
rect 934 3782 946 3834
rect 998 3782 1010 3834
rect 1062 3782 1080 3834
rect 664 3188 716 3194
rect 664 3130 716 3136
rect 800 2746 1080 3782
rect 1228 3777 1256 3878
rect 1214 3768 1270 3777
rect 1320 3754 1348 4542
rect 1412 3890 1440 4678
rect 2680 4378 2960 4400
rect 2680 4326 2698 4378
rect 2750 4326 2762 4378
rect 2814 4326 2826 4378
rect 2878 4326 2890 4378
rect 2942 4326 2960 4378
rect 1412 3862 1532 3890
rect 1320 3738 1440 3754
rect 1320 3732 1452 3738
rect 1320 3726 1400 3732
rect 1214 3703 1270 3712
rect 1400 3674 1452 3680
rect 1504 3670 1532 3862
rect 1492 3664 1544 3670
rect 1492 3606 1544 3612
rect 2680 3516 2960 4326
rect 2680 3460 2712 3516
rect 2768 3460 2792 3516
rect 2848 3460 2872 3516
rect 2928 3460 2960 3516
rect 2680 3436 2960 3460
rect 2680 3380 2712 3436
rect 2768 3380 2792 3436
rect 2848 3380 2872 3436
rect 2928 3380 2960 3436
rect 2680 3356 2960 3380
rect 2680 3300 2712 3356
rect 2768 3300 2792 3356
rect 2848 3300 2872 3356
rect 2928 3300 2960 3356
rect 2680 3290 2960 3300
rect 2680 3238 2698 3290
rect 2750 3238 2762 3290
rect 2814 3238 2826 3290
rect 2878 3238 2890 3290
rect 2942 3238 2960 3290
rect 1122 2952 1178 2961
rect 1122 2887 1124 2896
rect 1176 2887 1178 2896
rect 1124 2858 1176 2864
rect 800 2694 818 2746
rect 870 2694 882 2746
rect 934 2694 946 2746
rect 998 2694 1010 2746
rect 1062 2694 1080 2746
rect 800 2036 1080 2694
rect 1122 2680 1178 2689
rect 1122 2615 1124 2624
rect 1176 2615 1178 2624
rect 1124 2586 1176 2592
rect 1122 2408 1178 2417
rect 1122 2343 1178 2352
rect 800 1980 832 2036
rect 888 1980 912 2036
rect 968 1980 992 2036
rect 1048 1980 1080 2036
rect 800 1956 1080 1980
rect 1136 1970 1164 2343
rect 2680 2202 2960 3238
rect 2680 2150 2698 2202
rect 2750 2150 2762 2202
rect 2814 2150 2826 2202
rect 2878 2150 2890 2202
rect 2942 2150 2960 2202
rect 800 1900 832 1956
rect 888 1900 912 1956
rect 968 1900 992 1956
rect 1048 1900 1080 1956
rect 1124 1964 1176 1970
rect 1124 1906 1176 1912
rect 1308 1964 1360 1970
rect 1308 1906 1360 1912
rect 800 1876 1080 1900
rect 572 1828 624 1834
rect 572 1770 624 1776
rect 800 1820 832 1876
rect 888 1820 912 1876
rect 968 1820 992 1876
rect 1048 1820 1080 1876
rect 584 490 612 1770
rect 800 1658 1080 1820
rect 800 1606 818 1658
rect 870 1606 882 1658
rect 934 1606 946 1658
rect 998 1606 1010 1658
rect 1062 1606 1080 1658
rect 664 1420 716 1426
rect 664 1362 716 1368
rect 676 1193 704 1362
rect 662 1184 718 1193
rect 662 1119 718 1128
rect 800 1040 1080 1606
rect 1214 1592 1270 1601
rect 1214 1527 1216 1536
rect 1268 1527 1270 1536
rect 1216 1498 1268 1504
rect 1124 1488 1176 1494
rect 1124 1329 1176 1436
rect 1122 1320 1178 1329
rect 1122 1255 1178 1264
rect 754 490 810 600
rect 584 462 810 490
rect 754 -600 810 462
rect 1122 490 1178 600
rect 1320 490 1348 1906
rect 2680 1114 2960 2150
rect 2680 1062 2698 1114
rect 2750 1062 2762 1114
rect 2814 1062 2826 1114
rect 2878 1062 2890 1114
rect 2942 1062 2960 1114
rect 2680 1040 2960 1062
rect 1122 462 1348 490
rect 1122 -600 1178 462
<< via2 >>
rect 662 4392 718 4448
rect 1122 4004 1178 4040
rect 1122 3984 1124 4004
rect 1124 3984 1176 4004
rect 1176 3984 1178 4004
rect 1214 3712 1270 3768
rect 2712 3460 2768 3516
rect 2792 3460 2848 3516
rect 2872 3460 2928 3516
rect 2712 3380 2768 3436
rect 2792 3380 2848 3436
rect 2872 3380 2928 3436
rect 2712 3300 2768 3356
rect 2792 3300 2848 3356
rect 2872 3300 2928 3356
rect 1122 2916 1178 2952
rect 1122 2896 1124 2916
rect 1124 2896 1176 2916
rect 1176 2896 1178 2916
rect 1122 2644 1178 2680
rect 1122 2624 1124 2644
rect 1124 2624 1176 2644
rect 1176 2624 1178 2644
rect 1122 2352 1178 2408
rect 832 1980 888 2036
rect 912 1980 968 2036
rect 992 1980 1048 2036
rect 832 1900 888 1956
rect 912 1900 968 1956
rect 992 1900 1048 1956
rect 832 1820 888 1876
rect 912 1820 968 1876
rect 992 1820 1048 1876
rect 662 1128 718 1184
rect 1214 1556 1270 1592
rect 1214 1536 1216 1556
rect 1216 1536 1268 1556
rect 1268 1536 1270 1556
rect 1122 1264 1178 1320
<< metal3 >>
rect 657 4450 723 4453
rect 657 4448 858 4450
rect 657 4392 662 4448
rect 718 4392 858 4448
rect 657 4390 858 4392
rect 657 4387 723 4390
rect -600 4314 600 4344
rect 798 4314 858 4390
rect -600 4254 858 4314
rect -600 4224 600 4254
rect -600 4042 600 4072
rect 1117 4042 1183 4045
rect -600 4040 1183 4042
rect -600 3984 1122 4040
rect 1178 3984 1183 4040
rect -600 3982 1183 3984
rect -600 3952 600 3982
rect 1117 3979 1183 3982
rect -600 3770 600 3800
rect 1209 3770 1275 3773
rect -600 3768 1275 3770
rect -600 3712 1214 3768
rect 1270 3712 1275 3768
rect -600 3710 1275 3712
rect -600 3680 600 3710
rect 1209 3707 1275 3710
rect 412 3516 3268 3548
rect 412 3460 2712 3516
rect 2768 3460 2792 3516
rect 2848 3460 2872 3516
rect 2928 3460 3268 3516
rect 412 3436 3268 3460
rect 412 3380 2712 3436
rect 2768 3380 2792 3436
rect 2848 3380 2872 3436
rect 2928 3380 3268 3436
rect 412 3356 3268 3380
rect 412 3300 2712 3356
rect 2768 3300 2792 3356
rect 2848 3300 2872 3356
rect 2928 3300 3268 3356
rect 412 3268 3268 3300
rect -600 2954 600 2984
rect 1117 2954 1183 2957
rect -600 2952 1183 2954
rect -600 2896 1122 2952
rect 1178 2896 1183 2952
rect -600 2894 1183 2896
rect -600 2864 600 2894
rect 1117 2891 1183 2894
rect -600 2682 600 2712
rect 1117 2682 1183 2685
rect -600 2680 1183 2682
rect -600 2624 1122 2680
rect 1178 2624 1183 2680
rect -600 2622 1183 2624
rect -600 2592 600 2622
rect 1117 2619 1183 2622
rect -600 2410 600 2440
rect 1117 2410 1183 2413
rect -600 2408 1183 2410
rect -600 2352 1122 2408
rect 1178 2352 1183 2408
rect -600 2350 1183 2352
rect -600 2320 600 2350
rect 1117 2347 1183 2350
rect 412 2036 3268 2068
rect 412 1980 832 2036
rect 888 1980 912 2036
rect 968 1980 992 2036
rect 1048 1980 3268 2036
rect 412 1956 3268 1980
rect 412 1900 832 1956
rect 888 1900 912 1956
rect 968 1900 992 1956
rect 1048 1900 3268 1956
rect 412 1876 3268 1900
rect 412 1820 832 1876
rect 888 1820 912 1876
rect 968 1820 992 1876
rect 1048 1820 3268 1876
rect 412 1788 3268 1820
rect -600 1594 600 1624
rect 1209 1594 1275 1597
rect -600 1592 1275 1594
rect -600 1536 1214 1592
rect 1270 1536 1275 1592
rect -600 1534 1275 1536
rect -600 1504 600 1534
rect 1209 1531 1275 1534
rect -600 1322 600 1352
rect 1117 1322 1183 1325
rect -600 1320 1183 1322
rect -600 1264 1122 1320
rect 1178 1264 1183 1320
rect -600 1262 1183 1264
rect -600 1232 600 1262
rect 1117 1259 1183 1262
rect 657 1186 723 1189
rect 657 1184 858 1186
rect 657 1128 662 1184
rect 718 1128 858 1184
rect 657 1126 858 1128
rect 657 1123 723 1126
rect -600 1050 600 1080
rect 798 1050 858 1126
rect -600 990 858 1050
rect -600 960 600 990
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 1196 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1681316767
transform 1 0 1840 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18
timestamp 1681316767
transform 1 0 2116 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1681316767
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 736 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1681316767
transform 1 0 1288 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 1656 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1681316767
transform 1 0 2024 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_24
timestamp 1681316767
transform 1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1681316767
transform 1 0 736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 1288 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1681316767
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_26
timestamp 1681316767
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1681316767
transform 1 0 736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1681316767
transform 1 0 1288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_16
timestamp 1681316767
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp 1681316767
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1681316767
transform 1 0 736 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp 1681316767
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1681316767
transform 1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1681316767
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1681316767
transform 1 0 736 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_8
timestamp 1681316767
transform 1 0 1196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1681316767
transform 1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_18
timestamp 1681316767
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1681316767
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform -1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[1\]
timestamp 1681316767
transform -1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[2\]
timestamp 1681316767
transform -1 0 1196 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[3\]
timestamp 1681316767
transform -1 0 1840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[4\]
timestamp 1681316767
transform -1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[5\]
timestamp 1681316767
transform -1 0 1288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[6\]
timestamp 1681316767
transform -1 0 1288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[7\]
timestamp 1681316767
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[8\]
timestamp 1681316767
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[9\]
timestamp 1681316767
transform -1 0 1196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[10\]
timestamp 1681316767
transform -1 0 1288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[11\]
timestamp 1681316767
transform -1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  gpio_default_value\[12\]
timestamp 1681316767
transform -1 0 2024 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1681316767
transform 1 0 460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1681316767
transform -1 0 3220 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1681316767
transform 1 0 460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1681316767
transform -1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1681316767
transform 1 0 460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1681316767
transform -1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1681316767
transform 1 0 460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1681316767
transform -1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1681316767
transform 1 0 460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1681316767
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1681316767
transform 1 0 460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1681316767
transform -1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1681316767
transform 1 0 2024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1681316767
transform 1 0 2024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1681316767
transform 1 0 2024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1681316767
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
<< labels >>
flabel metal2 s 2680 1040 2960 4400 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 412 3268 3268 3548 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 800 1040 1080 4400 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 412 1788 3268 2068 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 754 5000 810 6200 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 2 nsew signal tristate
flabel metal3 s -600 4224 600 4344 0 FreeSans 480 0 0 0 gpio_defaults[10]
port 3 nsew signal tristate
flabel metal2 s 754 -600 810 600 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 4 nsew signal tristate
flabel metal2 s 1122 -600 1178 600 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 5 nsew signal tristate
flabel metal2 s 1122 5000 1178 6200 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 6 nsew signal tristate
flabel metal3 s -600 960 600 1080 0 FreeSans 480 0 0 0 gpio_defaults[2]
port 7 nsew signal tristate
flabel metal3 s -600 1232 600 1352 0 FreeSans 480 0 0 0 gpio_defaults[3]
port 8 nsew signal tristate
flabel metal3 s -600 1504 600 1624 0 FreeSans 480 0 0 0 gpio_defaults[4]
port 9 nsew signal tristate
flabel metal3 s -600 2320 600 2440 0 FreeSans 480 0 0 0 gpio_defaults[5]
port 10 nsew signal tristate
flabel metal3 s -600 2592 600 2712 0 FreeSans 480 0 0 0 gpio_defaults[6]
port 11 nsew signal tristate
flabel metal3 s -600 2864 600 2984 0 FreeSans 480 0 0 0 gpio_defaults[7]
port 12 nsew signal tristate
flabel metal3 s -600 3680 600 3800 0 FreeSans 480 0 0 0 gpio_defaults[8]
port 13 nsew signal tristate
flabel metal3 s -600 3952 600 4072 0 FreeSans 480 0 0 0 gpio_defaults[9]
port 14 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 3400 5600
<< end >>
